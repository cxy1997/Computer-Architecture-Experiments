`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:13:18 03/08/2017 
// Design Name: 
// Module Name:    Ledt_shift_2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Left_shift_2(INPUT, OUTPUT);
    input [31:0] INPUT;
	 output [31:0] OUTPUT;
	 assign OUTPUT = INPUT;

endmodule
