`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:49:41 03/27/2017 
// Design Name: 
// Module Name:    leftshift2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Left_shift_2(INPUT, OUTPUT);
    input [31:0] INPUT;
	 output [31:0] OUTPUT;
	 assign OUTPUT = INPUT;

endmodule